localparam N_GPIOS = 23;

localparam PIN_LED        = 0;

localparam PIN_DPAD_U     = 1;
localparam PIN_DPAD_D     = 2;
localparam PIN_DPAD_L     = 3;
localparam PIN_DPAD_R     = 4;
localparam PIN_BTN_A      = 5;
localparam PIN_BTN_B      = 6;
localparam PIN_BTN_X      = 7;
localparam PIN_BTN_Y      = 8;
localparam PIN_BTN_START  = 9;
localparam PIN_BTN_SELECT = 10;

localparam PIN_FLASH_CS   = 11;
localparam PIN_FLASH_SCLK = 12;
localparam PIN_FLASH_MOSI = 13;
localparam PIN_FLASH_MISO = 14;

localparam PIN_LCD_SCL    = 15;
localparam PIN_LCD_SDO    = 16;
localparam PIN_LCD_CS     = 17;
localparam PIN_LCD_DC     = 18;
localparam PIN_LCD_PWM    = 19;
localparam PIN_LCD_RST    = 20;

localparam PIN_UART_RX    = 21;
localparam PIN_UART_TX    = 22;
