always assume(rst_n == !$initstate);
always assume(!d_invalid);

always @ (posedge clk) begin

end