/******************************************************************************
 *     DO WHAT THE FUCK YOU WANT TO AND DON'T BLAME US PUBLIC LICENSE         *
 *                        Version 3, April 2008                               *
 *                                                                            *
 *     Copyright (C) 2019 Luke Wren                                           *
 *                                                                            *
 *     Everyone is permitted to copy and distribute verbatim or modified      *
 *     copies of this license document and accompanying software, and         *
 *     changing either is allowed.                                            *
 *                                                                            *
 *       TERMS AND CONDITIONS FOR COPYING, DISTRIBUTION AND MODIFICATION      *
 *                                                                            *
 *     0. You just DO WHAT THE FUCK YOU WANT TO.                              *
 *     1. We're NOT RESPONSIBLE WHEN IT DOESN'T FUCKING WORK.                 *
 *                                                                            *
 *****************************************************************************/

module hazard5_decode #(
	parameter EXTENSION_C = 1,   // compressed instruction extension
	parameter HAVE_CSR = 0,
	parameter W_ADDR = 32,
	parameter W_DATA = 32,
	parameter RESET_VECTOR = 32'h0,
	parameter W_REGADDR = 5
) (
	input wire clk,
	input wire rst_n,

	input wire  [31:0]          fd_cir,
	input wire  [1:0]           fd_cir_vld,
	output wire [1:0]           df_cir_use,
	output wire                 df_cir_lock,
	output reg                  d_jump_req,
	output reg  [W_ADDR-1:0]    d_jump_target,
	output wire [W_ADDR-1:0]    d_pc, // FIXME only added for riscv-formal

	output wire                 d_stall,
	input wire                  x_stall,
	input wire                  flush_d_x,
	input wire                  f_jump_rdy,
	input wire                  f_jump_now,
	input wire  [W_ADDR-1:0]    f_jump_target,

	output reg  [W_REGADDR-1:0] d_rs1, // combinatorial
	output reg  [W_REGADDR-1:0] d_rs2, // combinatorial

	output reg  [W_DATA-1:0]    dx_imm,
	output reg  [W_REGADDR-1:0] dx_rs1,
	output reg  [W_REGADDR-1:0] dx_rs2,
	output reg  [W_REGADDR-1:0] dx_rd,
	output reg  [W_ALUSRC-1:0]  dx_alusrc_a,
	output reg  [W_ALUSRC-1:0]  dx_alusrc_b,
	output reg  [W_ALUOP-1:0]   dx_aluop,
	output reg  [W_MEMOP-1:0]   dx_memop,
	output reg                  dx_csr_ren,
	output reg                  dx_csr_wen,
	output reg  [1:0]           dx_csr_wtype,
	output reg                  dx_csr_w_imm,
	output reg  [W_BCOND-1:0]   dx_branchcond,
	output reg  [W_ADDR-1:0]    dx_jump_target,
	output reg                  dx_jump_is_regoffs,
	output reg                  dx_result_is_linkaddr,
	output reg  [W_ADDR-1:0]    dx_pc,
	output reg  [W_ADDR-1:0]    dx_mispredict_addr,
	output reg  [2:0]           dx_except
);


// TODO TODO factor this out in a cleaner way, e.g. separate out registers and stall logic.

`include "rv_opcodes.vh"
`include "hazard5_ops.vh"

// ============================================================================
// PC/CIR control
// ============================================================================

wire d_starved = ~|fd_cir_vld || fd_cir_vld[0] && d_instr_is_32bit;
assign d_stall = x_stall ||
	d_starved || (d_jump_req && !f_jump_rdy);
assign df_cir_use =
	d_starved || d_stall ? 2'h0 :
	d_instr_is_32bit ? 2'h2 : 2'h1;

// CIR Locking is required if we successfully assert a jump request, but decode is stalled.
// (This only happens if decode stall is caused by X stall, not if fetch is starved!)
// The reason for this is that, if the CIR is not locked in, it can be trashed by
// incoming fetch data before the roadblock clears ahead of us, which will squash any other
// side effects this instruction may have besides jumping! This includes:
// - Linking for JAL
// - Mispredict recovery for branches
// Note that it is not possible to simply gate the jump request based on X stalling,
// because X stall is a function of hready, and jump request feeds haddr htrans etc.


wire assert_cir_lock = d_jump_req && f_jump_rdy && d_stall;
wire deassert_cir_lock = !d_stall;
reg cir_lock_prev;

assign df_cir_lock = (cir_lock_prev && !deassert_cir_lock) || assert_cir_lock;

always @ (posedge clk or negedge rst_n)
	if (!rst_n)
		cir_lock_prev <= 1'b0;
	else
		cir_lock_prev <= df_cir_lock;

reg  [W_ADDR-1:0]    pc;
wire [W_ADDR-1:0]    pc_next = pc + (d_instr_is_32bit ? 32'h4 : 32'h2);
assign d_pc = pc;

always @ (posedge clk or negedge rst_n) begin
	if (!rst_n) begin
		pc <= RESET_VECTOR;
	end else begin
		if ((f_jump_now && !assert_cir_lock) || (cir_lock_prev && deassert_cir_lock))
			pc <= f_jump_target;
		else if (!d_stall && !df_cir_lock)
			pc <= pc_next;
	end
end

// If the current CIR is there due to locking, it is a jump which has already had primary effect.
wire d_invalid;
wire jump_enable = !d_starved && !cir_lock_prev && !d_invalid;
reg [W_ADDR-1:0] d_jump_offs;


always @ (*) begin
	// JAL is major opcode 1101111,
	// branches are        1100011.
	case (d_instr[3])
	1'b1:    d_jump_offs = d_imm_j;
	default: d_jump_offs = d_imm_b;
	endcase

	d_jump_target = pc + d_jump_offs;

	casez ({d_instr[31], d_instr})
	{1'b1, RV_BEQ }: d_jump_req = jump_enable;
	{1'b1, RV_BNE }: d_jump_req = jump_enable;
	{1'b1, RV_BLT }: d_jump_req = jump_enable;
	{1'b1, RV_BGE }: d_jump_req = jump_enable;
	{1'b1, RV_BLTU}: d_jump_req = jump_enable;
	{1'b1, RV_BGEU}: d_jump_req = jump_enable;
	{1'bz, RV_JAL }: d_jump_req = jump_enable;
	default: d_jump_req = 1'b0;
	endcase
end

// ============================================================================
// Expand compressed instructions
// ============================================================================

wire [31:0] d_instr;
wire        d_instr_is_32bit;
wire        d_invalid_16bit;
reg         d_invalid_32bit;
assign      d_invalid = d_invalid_16bit || d_invalid_32bit;

hazard5_instr_decompress #(
	.PASSTHROUGH(!EXTENSION_C)
) decomp (
	.instr_in       (fd_cir),
	.instr_is_32bit (d_instr_is_32bit),
	.instr_out      (d_instr),
	.invalid        (d_invalid_16bit)
);

// ============================================================================
// Decode X controls
// ============================================================================

// Decode various immmediate formats
wire [31:0] d_imm_i = {{21{d_instr[31]}}, d_instr[30:20]};
wire [31:0] d_imm_s = {{21{d_instr[31]}}, d_instr[30:25], d_instr[11:7]};
wire [31:0] d_imm_b = {{20{d_instr[31]}}, d_instr[7], d_instr[30:25], d_instr[11:8], 1'b0};
wire [31:0] d_imm_u = {d_instr[31:12], {12{1'b0}}};
wire [31:0] d_imm_j = {{12{d_instr[31]}}, d_instr[19:12], d_instr[20], d_instr[30:21], 1'b0};

// Combinatorials:
reg  [W_REGADDR-1:0] d_rd;
reg  [W_DATA-1:0]    d_imm;
reg  [W_DATA-1:0]    d_branchoffs;
reg  [W_ALUSRC-1:0]  d_alusrc_a;
reg  [W_ALUSRC-1:0]  d_alusrc_b;
reg  [W_ALUOP-1:0]   d_aluop;
reg  [W_MEMOP-1:0]   d_memop;
reg  [W_BCOND-1:0]   d_branchcond;
reg                  d_jump_is_regoffs;
reg                  d_result_is_linkaddr;
reg                  d_csr_ren;
reg                  d_csr_wen;
reg  [1:0]           d_csr_wtype;
reg                  d_csr_w_imm;
reg  [W_EXCEPT-1:0]  d_except;

localparam X0 = {W_REGADDR{1'b0}};

always @ (*) begin
	// Assign some defaults
	d_rs1 = d_instr[19:15];
	d_rs2 = d_instr[24:20];
	d_rd  = d_instr[11: 7];
	d_imm = d_imm_i;
	d_branchoffs = d_imm_i;
	d_alusrc_a = ALUSRCA_RS1;
	d_alusrc_b = ALUSRCB_RS2;
	d_aluop = ALUOP_ADD;
	d_memop = MEMOP_NONE;
	d_csr_ren = 1'b0;
	d_csr_wen = 1'b0;
	d_csr_wtype = CSR_WTYPE_W;
	d_csr_w_imm = 1'b0;
	d_branchcond = BCOND_NEVER;
	d_jump_is_regoffs = 1'b0;
	d_result_is_linkaddr = 1'b0;
	d_invalid_32bit = 1'b0;
	d_except = EXCEPT_NONE;

	casez (d_instr)
	RV_BEQ:     begin d_rd = X0; d_aluop = ALUOP_SUB; d_branchcond = BCOND_ZERO;  end
	RV_BNE:     begin d_rd = X0; d_aluop = ALUOP_SUB; d_branchcond = BCOND_NZERO; end
	RV_BLT:     begin d_rd = X0; d_aluop = ALUOP_LT;  d_branchcond = BCOND_NZERO; end
	RV_BGE:     begin d_rd = X0; d_aluop = ALUOP_LT;  d_branchcond = BCOND_ZERO; end
	RV_BLTU:    begin d_rd = X0; d_aluop = ALUOP_LTU; d_branchcond = BCOND_NZERO; end
	RV_BGEU:    begin d_rd = X0; d_aluop = ALUOP_LTU; d_branchcond = BCOND_ZERO; end
	RV_JALR:    begin d_result_is_linkaddr = 1'b1; d_jump_is_regoffs = 1'b1; d_aluop = ALUOP_ADD; d_imm = d_imm_i; d_alusrc_b = ALUSRCB_IMM; d_rs2 = X0; d_branchcond = BCOND_ALWAYS; end
	RV_JAL:     begin d_result_is_linkaddr = 1'b1; d_rs2 = X0; d_rs1 = X0; end
	RV_LUI:     begin d_aluop = ALUOP_ADD; d_imm = d_imm_u; d_alusrc_b = ALUSRCB_IMM; d_rs2 = X0; d_rs1 = X0; end
	RV_AUIPC:   begin d_aluop = ALUOP_ADD; d_imm = d_imm_u; d_alusrc_b = ALUSRCB_IMM; d_rs2 = X0; d_alusrc_a = ALUSRCA_PC;  d_rs1 = X0; end
	RV_ADDI:    begin d_aluop = ALUOP_ADD; d_imm = d_imm_i; d_alusrc_b = ALUSRCB_IMM; d_rs2 = X0; end
	RV_SLLI:    begin d_aluop = ALUOP_SLL; d_imm = d_imm_i; d_alusrc_b = ALUSRCB_IMM; d_rs2 = X0; end
	RV_SLTI:    begin d_aluop = ALUOP_LT;  d_imm = d_imm_i; d_alusrc_b = ALUSRCB_IMM; d_rs2 = X0; end
	RV_SLTIU:   begin d_aluop = ALUOP_LTU; d_imm = d_imm_i; d_alusrc_b = ALUSRCB_IMM; d_rs2 = X0; end
	RV_XORI:    begin d_aluop = ALUOP_XOR; d_imm = d_imm_i; d_alusrc_b = ALUSRCB_IMM; d_rs2 = X0; end
	RV_SRLI:    begin d_aluop = ALUOP_SRL; d_imm = d_imm_i; d_alusrc_b = ALUSRCB_IMM; d_rs2 = X0; end
	RV_SRAI:    begin d_aluop = ALUOP_SRA; d_imm = d_imm_i; d_alusrc_b = ALUSRCB_IMM; d_rs2 = X0; end
	RV_ORI:     begin d_aluop = ALUOP_OR;  d_imm = d_imm_i; d_alusrc_b = ALUSRCB_IMM; d_rs2 = X0; end
	RV_ANDI:    begin d_aluop = ALUOP_AND; d_imm = d_imm_i; d_alusrc_b = ALUSRCB_IMM; d_rs2 = X0; end
	RV_ADD:     begin d_aluop = ALUOP_ADD; end
	RV_SUB:     begin d_aluop = ALUOP_SUB; end
	RV_SLL:     begin d_aluop = ALUOP_SLL; end
	RV_SLT:     begin d_aluop = ALUOP_LT;  end
	RV_SLTU:    begin d_aluop = ALUOP_LTU; end
	RV_XOR:     begin d_aluop = ALUOP_XOR; end
	RV_SRL:     begin d_aluop = ALUOP_SRL; end
	RV_SRA:     begin d_aluop = ALUOP_SRA; end
	RV_OR:      begin d_aluop = ALUOP_OR;  end
	RV_AND:     begin d_aluop = ALUOP_AND; end
	RV_LB:      begin d_aluop = ALUOP_ADD; d_imm = d_imm_i; d_alusrc_b = ALUSRCB_IMM; d_rs2 = X0; d_memop = MEMOP_LB;  end
	RV_LH:      begin d_aluop = ALUOP_ADD; d_imm = d_imm_i; d_alusrc_b = ALUSRCB_IMM; d_rs2 = X0; d_memop = MEMOP_LH;  end
	RV_LW:      begin d_aluop = ALUOP_ADD; d_imm = d_imm_i; d_alusrc_b = ALUSRCB_IMM; d_rs2 = X0; d_memop = MEMOP_LW;  end
	RV_LBU:     begin d_aluop = ALUOP_ADD; d_imm = d_imm_i; d_alusrc_b = ALUSRCB_IMM; d_rs2 = X0; d_memop = MEMOP_LBU; end
	RV_LHU:     begin d_aluop = ALUOP_ADD; d_imm = d_imm_i; d_alusrc_b = ALUSRCB_IMM; d_rs2 = X0; d_memop = MEMOP_LHU; end
	RV_SB:      begin d_aluop = ALUOP_ADD; d_imm = d_imm_s; d_alusrc_b = ALUSRCB_IMM; d_memop = MEMOP_SB;  d_rd = X0; end
	RV_SH:      begin d_aluop = ALUOP_ADD; d_imm = d_imm_s; d_alusrc_b = ALUSRCB_IMM; d_memop = MEMOP_SH;  d_rd = X0; end
	RV_SW:      begin d_aluop = ALUOP_ADD; d_imm = d_imm_s; d_alusrc_b = ALUSRCB_IMM; d_memop = MEMOP_SW;  d_rd = X0; end
	RV_FENCE:   begin d_rd = X0; end  // NOP
	RV_FENCE_I: begin d_rd = X0; end  // NOP // TODO: this should be jump to PC + 4. Evaluate the cost of doing this in decode (or find a way of doing it in X).
	RV_CSRRW:   if (HAVE_CSR) begin d_imm = d_imm_i; d_csr_wen = 1'b1  ; d_csr_ren = |d_rd; d_csr_wtype = CSR_WTYPE_W; end else begin d_invalid_32bit = 1'b1; end
	RV_CSRRS:   if (HAVE_CSR) begin d_imm = d_imm_i; d_csr_wen = |d_rs1; d_csr_ren = 1'b1 ; d_csr_wtype = CSR_WTYPE_S; end else begin d_invalid_32bit = 1'b1; end
	RV_CSRRC:   if (HAVE_CSR) begin d_imm = d_imm_i; d_csr_wen = |d_rs1; d_csr_ren = 1'b1 ; d_csr_wtype = CSR_WTYPE_C; end else begin d_invalid_32bit = 1'b1; end
	RV_CSRRWI:  if (HAVE_CSR) begin d_imm = d_imm_i; d_csr_wen = 1'b1  ; d_csr_ren = |d_rd; d_csr_wtype = CSR_WTYPE_W; d_csr_w_imm = 1'b1; end else begin d_invalid_32bit = 1'b1; end
	RV_CSRRSI:  if (HAVE_CSR) begin d_imm = d_imm_i; d_csr_wen = |d_rs1; d_csr_ren = 1'b1 ; d_csr_wtype = CSR_WTYPE_S; d_csr_w_imm = 1'b1; end else begin d_invalid_32bit = 1'b1; end
	RV_CSRRCI:  if (HAVE_CSR) begin d_imm = d_imm_i; d_csr_wen = |d_rs1; d_csr_ren = 1'b1 ; d_csr_wtype = CSR_WTYPE_C; d_csr_w_imm = 1'b1; end else begin d_invalid_32bit = 1'b1; end
	RV_ECALL:   begin d_except = EXCEPT_ECALL;  d_rs2 = X0; d_rs1 = X0; d_rd = X0; end
	RV_EBREAK:  begin d_except = EXCEPT_EBREAK; d_rs2 = X0; d_rs1 = X0; d_rd = X0; end
	RV_MRET:    begin d_except = EXCEPT_MRET;   d_rs2 = X0; d_rs1 = X0; d_rd = X0; end
	RV_SYSTEM:  begin
		//synthesis translate_off
		if (!d_stall && !clk) $display("Syscall @ PC %h: %h", pc, d_instr);
		//synthesis translate_on
		d_except = EXCEPT_INSTR_ILLEGAL; d_rs2 = X0; d_rs1 = X0; d_rd = X0;
	 end
	default:    begin d_invalid_32bit = 1'b1; end
	endcase
end


always @ (posedge clk or negedge rst_n) begin
	if (!rst_n) begin
		{dx_rs1, dx_rs2, dx_rd} <= {(3 * W_REGADDR){1'b0}};
		dx_alusrc_a <= ALUSRCA_RS1;
		dx_alusrc_b <= ALUSRCB_RS2;
		dx_aluop <= ALUOP_ADD;
		dx_memop <= MEMOP_NONE;
		dx_csr_ren <= 1'b0;
		dx_csr_wen <= 1'b0;
		dx_csr_wtype <= CSR_WTYPE_W;
		dx_csr_w_imm <= 1'b0;
		dx_branchcond <= BCOND_NEVER;
		dx_jump_is_regoffs <= 1'b0;
		dx_result_is_linkaddr <= 1'b0;
		dx_except <= EXCEPT_NONE;
	end else if (!x_stall) begin
		// These ones can have side effects
		dx_rs1        <= d_invalid ? {W_REGADDR{1'b0}}    : d_rs1;
		dx_rs2        <= d_invalid ? {W_REGADDR{1'b0}}    : d_rs2;
		dx_rd         <= d_invalid ? {W_REGADDR{1'b0}}    : d_rd;
		dx_memop      <= d_invalid ? MEMOP_NONE           : d_memop;
		dx_branchcond <= d_invalid ? BCOND_NEVER          : d_branchcond;
		dx_csr_ren    <= d_invalid ? 1'b0                 : d_csr_ren;
		dx_csr_wen    <= d_invalid ? 1'b0                 : d_csr_wen;
		dx_except     <= d_invalid ? EXCEPT_INSTR_ILLEGAL : d_except;

		// These can't
		dx_alusrc_a <= d_alusrc_a;
		dx_alusrc_b <= d_alusrc_b;
		dx_aluop <= d_aluop;
		dx_jump_is_regoffs <= d_jump_is_regoffs;
		dx_result_is_linkaddr <= d_result_is_linkaddr;
		dx_csr_wtype <= d_csr_wtype;
		dx_csr_w_imm <= d_csr_w_imm;

		// Bubble insertion
		if (d_stall || flush_d_x) begin
			dx_branchcond <= BCOND_NEVER;
			dx_memop <= MEMOP_NONE;
			dx_rd <= 5'h0;
			dx_except <= EXCEPT_NONE;
			dx_csr_ren <= 1'b0;
			dx_csr_wen <= 1'b0;
			// Also need to clear rs1, rs2, due to a nasty sequence of events:
			// Suppose we have a load, followed by a dependent branch, which is predicted taken
			// - branch will stall in D until AHB master becomes free
			// - on next cycle, prediction causes jump, and bubble is in X
			// - if X gets branch's rs1, rs2, it will cause spurious RAW stall
			// - on next cycle, branch will not progress into X due to RAW stall, but *will* be replaced in D due to jump
			// - branch mispredict now cannot be corrected
			dx_rs1 <= 5'h0;
			dx_rs2 <= 5'h0;
		end
	end
end

// No reset required on these; will be masked by the resettable pipeline controls until they're valid
always @ (posedge clk) begin
	if (!x_stall) begin
		dx_imm <= d_imm;
		dx_jump_target <= d_jump_target;
		dx_pc <= pc;
		dx_mispredict_addr <= pc_next;
	end
end

endmodule
