localparam N_GPIOS = 11;

localparam PIN_LED        = 0;

localparam PIN_DPAD_U     = 1;
localparam PIN_DPAD_D     = 2;
localparam PIN_DPAD_L     = 3;
localparam PIN_DPAD_R     = 4;
localparam PIN_BTN_A      = 5;
localparam PIN_BTN_B      = 6;
localparam PIN_BTN_X      = 7;
localparam PIN_BTN_Y      = 8;
localparam PIN_BTN_START  = 9;
localparam PIN_BTN_SELECT = 10;
